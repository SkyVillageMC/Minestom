{"0,122,9":1,"14,122,8":1,"14,122,9":1,"0,122,7":1,"0,122,8":1,"14,122,4":1,"14,122,5":1,"14,122,6":1,"14,122,7":1,"6,122,0":1,"14,122,0":1,"14,122,1":1,"14,122,2":1,"14,122,3":1,"15,123,8":1,"7,124,6":1,"8,122,11":1,"8,122,10":1,"6,123,6":1,"6,123,5":1,"6,123,4":1,"4,122,12":1,"4,122,13":1,"4,122,14":1,"6,122,15":1,"4,122,15":1,"6,122,14":1,"6,122,13":1,"2,122,12":1,"6,122,12":1,"2,122,13":1,"6,122,11":1,"0,122,10":1,"2,122,10":1,"4,122,10":1,"4,122,11":1,"2,122,11":1,"0,122,11":1,"6,122,10":1,"5,124,12":1,"0,122,12":1,"8,122,13":1,"0,122,13":1,"8,122,12":1,"2,122,14":1,"0,122,14":1,"8,122,15":1,"2,122,15":1,"0,122,15":1,"8,122,14":1,"15,122,2":1,"15,122,1":1,"15,122,0":1,"15,122,6":1,"15,122,5":1,"15,122,4":1,"7,125,4":1,"15,122,3":1,"15,122,9":1,"15,122,8":1,"15,122,7":1,"13,123,13":1,"7,125,6":1,"7,125,5":1,"6,124,6":1,"6,124,5":1,"6,124,4":1,"12,122,15":1,"12,122,14":1,"12,122,13":1,"8,125,4":1,"8,125,5":1,"8,125,6":1,"12,122,12":1,"11,124,13":1,"12,122,11":1,"12,122,10":1,"5,123,9":1,"8,123,12":1,"10,122,3":1,"10,122,2":1,"10,122,1":1,"10,122,0":1,"10,122,7":1,"10,122,6":1,"10,122,5":1,"10,122,4":1,"7,122,5":1,"7,122,4":1,"3,123,13":1,"7,122,7":1,"10,122,9":1,"7,122,6":1,"10,122,8":1,"7,122,1":1,"5,123,12":1,"2,123,13":1,"7,122,0":1,"7,122,3":1,"0,123,11":1,"2,123,11":1,"7,122,2":1,"2,123,12":1,"3,123,11":1,"0,123,13":1,"0,123,14":1,"2,123,15":1,"7,122,9":1,"7,122,8":1,"4,122,6":1,"4,122,5":1,"4,122,4":1,"13,122,9":1,"4,122,3":1,"13,122,7":1,"4,122,9":1,"13,122,8":1,"4,122,8":1,"13,122,5":1,"4,122,7":1,"13,122,6":1,"13,122,14":1,"8,124,5":1,"13,122,15":1,"8,124,6":1,"5,122,1":1,"5,122,0":1,"13,122,3":1,"13,122,10":1,"15,122,15":1,"13,122,4":1,"13,122,11":1,"15,122,14":1,"13,122,1":1,"13,122,12":1,"15,122,13":1,"13,122,2":1,"13,122,13":1,"15,122,12":1,"8,124,4":1,"15,122,11":1,"13,122,0":1,"15,122,10":1,"12,122,6":1,"12,122,7":1,"12,122,8":1,"12,122,9":1,"5,122,3":1,"5,122,2":1,"5,122,5":1,"14,123,9":1,"5,122,4":1,"5,122,7":1,"5,122,6":1,"5,122,9":1,"5,122,8":1,"7,123,6":1,"12,123,11":1,"12,122,0":1,"12,122,1":1,"12,123,13":1,"15,123,13":1,"12,122,2":1,"12,122,3":1,"15,123,11":1,"12,122,4":1,"12,122,5":1,"11,122,1":1,"11,122,2":1,"11,122,0":1,"11,122,5":1,"11,122,6":1,"11,122,3":1,"6,122,9":1,"11,122,4":1,"6,122,8":1,"6,122,7":1,"6,122,6":1,"6,122,5":1,"6,122,4":1,"6,122,3":1,"6,122,2":1,"6,122,1":1,"3,122,10":1,"10,122,12":1,"10,122,11":1,"10,122,14":1,"10,122,13":1,"3,122,14":1,"8,123,6":1,"3,122,13":1,"10,122,15":1,"3,122,12":1,"3,122,11":1,"11,122,9":1,"11,122,7":1,"8,123,4":1,"3,122,15":1,"11,122,8":1,"8,123,5":1,"10,122,10":1,"3,122,1":1,"3,122,0":1,"3,122,3":1,"3,122,2":1,"8,122,7":1,"8,122,8":1,"8,122,9":1,"8,122,3":1,"3,123,8":1,"12,124,11":1,"8,122,4":1,"8,122,5":1,"8,122,6":1,"8,122,0":1,"8,122,1":1,"8,122,2":1,"2,122,9":1,"2,122,7":1,"2,122,8":1,"2,122,5":1,"2,122,6":1,"14,123,13":1,"4,122,2":1,"14,123,10":1,"4,122,1":1,"14,123,11":1,"4,122,0":1,"9,122,0":1,"9,122,1":1,"9,122,4":1,"9,122,11":1,"9,122,5":1,"9,122,12":1,"9,122,2":1,"9,122,3":1,"9,122,10":1,"9,122,8":1,"9,122,9":1,"9,122,6":1,"9,122,7":1,"5,122,14":1,"5,122,13":1,"5,122,15":1,"1,122,10":1,"5,122,10":1,"0,124,11":1,"1,122,12":1,"5,122,12":1,"1,122,11":1,"5,122,11":1,"1,122,14":1,"3,122,9":1,"9,122,15":1,"1,122,13":1,"3,122,8":1,"9,122,13":1,"1,122,15":1,"9,122,14":1,"3,122,5":1,"3,122,4":1,"3,122,7":1,"3,122,6":1,"9,123,12":1,"7,123,11":1,"1,123,11":1,"6,123,11":1,"7,123,12":1,"6,125,6":1,"2,122,3":1,"6,125,5":1,"2,122,4":1,"6,125,4":1,"2,122,1":1,"2,122,2":1,"2,122,0":1,"1,122,6":1,"11,122,14":1,"1,122,7":1,"11,122,15":1,"1,122,8":1,"11,122,12":1,"1,122,9":1,"11,122,13":1,"11,122,10":1,"11,122,11":1,"1,122,0":1,"1,122,1":1,"1,122,2":1,"1,122,3":1,"1,122,4":1,"1,122,5":1,"11,123,13":1,"11,123,12":1,"7,122,10":1,"0,122,1":1,"0,122,2":1,"1,123,7":1,"0,122,0":1,"0,122,5":1,"0,122,6":1,"14,122,15":1,"0,122,3":1,"0,122,4":1,"7,122,11":1,"14,122,12":1,"7,122,12":1,"14,122,11":1,"7,122,13":1,"14,122,14":1,"7,122,14":1,"14,122,13":1,"7,122,15":1,"14,122,10":1}